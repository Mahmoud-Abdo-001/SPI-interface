package fsm_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "fsm_sequence_item.sv"
    `include "fsm_monitor.sv"
    `include "fsm_agent.sv"
    `include "fsm_scoreboard.sv"
    `include "fsm_coverage_collector.sv"

endpackage