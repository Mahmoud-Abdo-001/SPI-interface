package ram_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ram_sequence_item.sv"
    `include "ram_monitor.sv"
    `include "ram_agent.sv"
    `include "ram_scoreboard.sv"
    `include "ram_coverage_collector.sv"

endpackage